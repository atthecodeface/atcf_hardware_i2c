/** Copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_apb_target_i2c.cdl
 * @brief Testbench for APB processor (ROM-based APB trasanctions)
 *
 * This is a simple testbench for the ROM-based APB transaction processor
 */
/*a Includes */
include "apb::apb.h"
include "apb::apb_targets.h"
include "i2c.h"
include "i2c_modules.h"

/*a Module */
module tb_apb_target_i2c( clock clk,
                          input bit reset_n,
                          input t_apb_request   apb_request,
                          output t_apb_response apb_response,
                          output t_i2c i2c_in,
                          input  t_i2c i2c_th,
                          input  t_i2c_conf i2c_conf,
                          output bit[16] gpio_output,
                          output bit[16] gpio_output_enable
)
{

    /*b Nets */
    comb t_apb_request[2]   apb_request_mod;
    net  t_apb_response[2]  apb_response_mod;
    net t_apb_request   i2c_apb_request;
    net t_apb_response  i2c_apb_response;
    net t_i2c i2c_slave;
    net t_i2c[2] i2c_master;

    comb t_i2c_slave_select slave_select;
    net t_i2c_action i2c_action;
    net t_i2c_slave_request slave_request;
    net t_i2c_slave_response slave_response;
    net bit[16] gpio_output;
    net bit[16] gpio_output_enable;

    /*b Instantiations */
    instantiations: {
        i2c_in  = i2c_th;
        // i2c_in &= i2c_slave;
        i2c_in.scl = i2c_in.scl & i2c_slave.scl;
        i2c_in.sda = i2c_in.sda & i2c_slave.sda;
        for (i; 2) {
            i2c_in.scl = i2c_in.scl & i2c_master[i].scl;
            i2c_in.sda = i2c_in.sda & i2c_master[i].sda;
        }
        slave_select = {mask=7h70, value=7h10};

        apb_response = {*=0};
        for (i; 2) {
            apb_request_mod[i]      = apb_request;
            apb_request_mod[i].psel = apb_request.psel && (apb_request.paddr[4;16]==i);
            apb_response           |= apb_response_mod[i];
        }
        for (i; 2) {
            apb_target_i2c_master apb_i2c[i]( clk <- clk,
                                              reset_n <= reset_n,
                                              apb_request  <= apb_request_mod[i],
                                              apb_response => apb_response_mod[i],
                                              i2c_in  <= i2c_in,
                                              i2c_out => i2c_master[i] );
        }

        i2c_interface i2c( clk <- clk,
                           reset_n <= reset_n,
                           i2c_in <= i2c_in,
                           i2c_action => i2c_action,
                           i2c_conf <= i2c_conf );
        
        i2c_slave slave(clk <- clk,
                        reset_n    <= reset_n,
                        i2c_action <= i2c_action,
                        i2c_out    => i2c_slave,
                        slave_select   <= slave_select, 
                        slave_request  => slave_request,
                        slave_response <= slave_response );

        i2c_slave_apb_master i2c_apb( clk <- clk,
                                      reset_n <= reset_n,
                                      slave_request <= slave_request,
                                      slave_response => slave_response,
                                      apb_request => i2c_apb_request,
                                      apb_response <= i2c_apb_response );
        apb_target_gpio gpio(clk <- clk,
                             reset_n <= reset_n,
                             apb_request <= i2c_apb_request,
                             apb_response => i2c_apb_response,
                             gpio_output => gpio_output,
                             gpio_output_enable => gpio_output_enable,
                             gpio_input <= gpio_output);
    }

    /*b All done */
}
